TOP/statementlist.0.9:
  statement/EXPR/value/number.1.3:
    integer/decint.1.3: null
  statement/EXPR/value/number.4.7:
    integer/VALUE.4.7: null
